//--------------------------------------------------------------------------------------------------
// Design    : nova
// Author(s) : Ke Xu
// Email	   : eexuke@yahoo.com
// File      : hybrid_pipeline_ctrl.v
// Generated : Sept 5, 2005
// Copyright (C) 2008 Ke Xu                
//-------------------------------------------------------------------------------------------------
// Description 
// Control 4x4 block level pipeline for reconstruction
// Receive the 1cycle end_of_xxx signal(combinational)
// Generated the 1cycle trigger_xxx signal
//-------------------------------------------------------------------------------------------------
// Revise log 
// 1.April 11,2006
// Modify the 1cycle trigger_xxx signal from registers to combinational logic to save decoding clock cycles
//-------------------------------------------------------------------------------------------------

// synopsys translate_off
//`include "timescale.v"
// synopsys translate_on
`include "nova_defines.v"

module hybrid_pipeline_ctrl (clk,reset_n,mb_num_h,mb_num_v,blk4x4_rec_counter,CodedBlockPatternLuma,CodedBlockPatternChroma,
	mb_type_general,slice_data_state,residual_state,TotalCoeff,Is_skip_run_entry,skip_mv_calc,
	end_of_one_residual_block,end_of_DCBlk_IQIT,end_of_ACBlk4x4_IQIT,end_of_one_blk4x4_intra,end_of_one_blk4x4_inter,
	end_of_one_blk4x4_sum,end_of_MB_DF,disable_DF,
	
	curr_CBPLuma_IsZero,end_of_MB_DEC,trigger_CAVLC,trigger_blk4x4_intra_pred,
	trigger_blk4x4_inter_pred,trigger_blk4x4_rec_sum);
	input clk,reset_n;
	input [3:0] mb_num_h;
	input [3:0] mb_num_v;
	input [4:0] blk4x4_rec_counter;
	input [3:0] CodedBlockPatternLuma;
	input [1:0] CodedBlockPatternChroma;
	input [3:0] mb_type_general;
	input [3:0] slice_data_state;
	input [3:0] residual_state;
	input [4:0] TotalCoeff;
	input Is_skip_run_entry;
	input skip_mv_calc;
	input end_of_one_residual_block;
	input end_of_DCBlk_IQIT;
	input end_of_ACBlk4x4_IQIT;
	input end_of_one_blk4x4_intra,end_of_one_blk4x4_inter,end_of_one_blk4x4_sum;
	input end_of_MB_DF;
	input disable_DF;
	
	output curr_CBPLuma_IsZero;
	output end_of_MB_DEC;
	output trigger_CAVLC;
	output trigger_blk4x4_intra_pred,trigger_blk4x4_inter_pred;
	output trigger_blk4x4_rec_sum;
	
	//change trigger_blk4x4_intra_pred from combination to reg
	reg trigger_CAVLC;             //combination
	reg trigger_blk4x4_intra_pred; //reg
	reg trigger_blk4x4_inter_pred; //reg
	reg trigger_blk4x4_rec_sum;    //combination
	
	//CBPLuma only make sense for residual_state == LumaLevel_s
	//CBPLuma is derived to help judge whether res_blk4x4_IsAllZero caused by CodedBlockPattern != 4'b1111
	reg curr_CBPLuma_IsZero;
	always @ (blk4x4_rec_counter or CodedBlockPatternLuma)
		if (blk4x4_rec_counter < 16)
			case (blk4x4_rec_counter[3:2])
				2'b00:curr_CBPLuma_IsZero <= !CodedBlockPatternLuma[0];
				2'b01:curr_CBPLuma_IsZero <= !CodedBlockPatternLuma[1];
				2'b10:curr_CBPLuma_IsZero <= !CodedBlockPatternLuma[2]; 
				2'b11:curr_CBPLuma_IsZero <= !CodedBlockPatternLuma[3];
			endcase
		else
			curr_CBPLuma_IsZero <= 0;
	//---------------------------------------------------------------------------------
	//signals to trigger:
	//	1.4x4 blk CAVLC
	//	2.4x4 Intra Prediction
	//	3.4x4 Inter Prediction 
	//	4.4x4 reconstruction sum
	//	5.16x16 deblocking filter
	//	All the trigger_xxx signals are generated by sequential logic
	//---------------------------------------------------------------------------------	
	
	//1. trigger_CAVLC: when reconstruction is dealing with skip_run or zero residual (construction 
	//   only from inter/intra prediction) blocks,CAVLC decoder,as well as whole bitstream parsing FSM,
	//   needs to be stalled and wait until the reconstruction process of previous 
 
	always @ (slice_data_state or residual_state or mb_type_general[3:2] or CodedBlockPatternLuma 
		or CodedBlockPatternChroma or end_of_one_residual_block or end_of_DCBlk_IQIT or end_of_one_blk4x4_sum 
		or blk4x4_rec_counter or TotalCoeff or curr_CBPLuma_IsZero)
		//	Entry
		if (slice_data_state == `residual && residual_state == `rst_residual)
			begin
				if (mb_type_general[3:2] == 2'b10)			//Intra16x16:first block must be DC
					trigger_CAVLC <= 1'b1;
				else if (CodedBlockPatternLuma[0] == 1'b0)	//First 8x8 block has no residuals
					trigger_CAVLC <= 1'b0;
				else  										//normal case
					trigger_CAVLC <= 1'b1;
			end	
		//	End of one DC
		else if ((residual_state == `Intra16x16DCLevel_s || residual_state == `ChromaDCLevel_Cb_s ||
		residual_state == `ChromaDCLevel_Cr_s) && ((end_of_one_residual_block && TotalCoeff == 0)|| end_of_DCBlk_IQIT))
			case (residual_state)
				`Intra16x16DCLevel_s:	//end of luma DC
				trigger_CAVLC <= (CodedBlockPatternLuma[0] == 1'b0)? 1'b0:1'b1;
				`ChromaDCLevel_Cb_s:		//end of chroma DC Cb,trigger chroma DC Cr now!
				trigger_CAVLC <= 1'b1;
				`ChromaDCLevel_Cr_s:		//end of chroma DC Cr
				trigger_CAVLC <= (CodedBlockPatternChroma == 2'b01)? 1'b0:1'b1;
				default:trigger_CAVLC <= 1'b0;
			endcase
		//	End of skip or normal
		else if (end_of_one_blk4x4_sum)
			begin
				if (slice_data_state == `skip_run_duration)
					trigger_CAVLC <= 1'b0;
				else 
					case (blk4x4_rec_counter)
						0,1,2,4,5,6,8,9,10,12,13,14:trigger_CAVLC <= (curr_CBPLuma_IsZero)? 1'b0:1'b1;
						3 :trigger_CAVLC <= (CodedBlockPatternLuma[1])? 1'b1:1'b0;
						7 :trigger_CAVLC <= (CodedBlockPatternLuma[2])? 1'b1:1'b0;
						11:trigger_CAVLC <= (CodedBlockPatternLuma[3])? 1'b1:1'b0;
						15:trigger_CAVLC <= (CodedBlockPatternChroma == 0)? 1'b0:1'b1;
						23:trigger_CAVLC <= 1'b0;
						default:trigger_CAVLC <= (CodedBlockPatternChroma == 2)? 1'b1:1'b0;
					endcase
			end
		else
			trigger_CAVLC <= 1'b0;
	
	//end_of_MB_rec:end of one MB reconstruction 
	wire end_of_MB_rec;
	assign end_of_MB_rec = (blk4x4_rec_counter == 5'd23 && end_of_one_blk4x4_sum == 1'b1)? 1'b1:1'b0;
	
	//MB_needs_DF: identify whether this MB needs to be deblocking filtered
	reg MB_needs_DF;
	always @ (posedge clk)
		if (reset_n == 1'b0)
			MB_needs_DF <= 1'b0;
		else if (end_of_MB_DEC == 1'b1 && !disable_DF)
			MB_needs_DF <= 1'b1;
		else if (end_of_MB_DEC == 1'b1 && disable_DF)
			MB_needs_DF <= 1'b0;
	//MB_rec_DF_align:latch the first arrival of end_of_MB_rec and end_of_MB_DF
	reg MB_rec_DF_align;
	always @ (posedge clk)
		if (reset_n == 1'b0)
			MB_rec_DF_align <= 1'b0;
		else if (end_of_MB_DEC)
			MB_rec_DF_align <= 1'b0;
		else if (MB_needs_DF && (end_of_MB_rec || end_of_MB_DF == 1'b1))
			MB_rec_DF_align <= 1'b1;
		 
			
	//end_of_MB_DEC:end of one macroblock decoding (end of both reconstruction and previous MB's deblocking
	// (if previous MB needs deblocking)),generated by combinational logic
	reg end_of_MB_DEC;
	always @ (MB_needs_DF or end_of_MB_rec or end_of_MB_DF or MB_rec_DF_align or mb_num_h or mb_num_v)
		if (MB_needs_DF == 1'b1)
			begin
				if (end_of_MB_rec && end_of_MB_DF)	//arrive simultaneously
					end_of_MB_DEC <= 1'b1;
				else if (MB_rec_DF_align == 1'b1 && (end_of_MB_rec || end_of_MB_DF))
					end_of_MB_DEC <= 1'b1;
				else if (mb_num_h == 0 && mb_num_v == 0 && end_of_MB_rec)//first MB has no correspinding DF process
					end_of_MB_DEC <= 1'b1;
				else
					end_of_MB_DEC <= 1'b0;
			end
		else
			end_of_MB_DEC <= (end_of_MB_rec)? 1'b1:1'b0;
			
	//2. trigger_blk4x4_intra_pred
	wire trigger_blk4x4_intra_pred_tmp;
	assign trigger_blk4x4_intra_pred_tmp = (mb_type_general[3] && ((slice_data_state == `residual && 
	residual_state == `rst_residual) || (end_of_one_blk4x4_sum && blk4x4_rec_counter != 23)))? 1'b1:1'b0;
	
	always @ (posedge clk)
		if (reset_n == 1'b0)
			trigger_blk4x4_intra_pred <= 1'b0;
		else
			trigger_blk4x4_intra_pred <= trigger_blk4x4_intra_pred_tmp;
			
	//3. trigger_blk4x4_inter_pred
	always @ (posedge clk)
		if (reset_n == 1'b0)
			trigger_blk4x4_inter_pred <= 1'b0;
		//For skip_run_duration
		// 1.trigger inter pred when entering skip_run_duration after mb_skip_run_s state
		else if (Is_skip_run_entry)
			trigger_blk4x4_inter_pred <= 1'b1;
		// 2.trigger inter pred during skip_run_duration
		else if (slice_data_state == `skip_run_duration)
			begin
				if (skip_mv_calc)
					trigger_blk4x4_inter_pred <= 1'b1;
				else 
					trigger_blk4x4_inter_pred <= (end_of_one_blk4x4_sum && blk4x4_rec_counter != 23)? 1'b1:1'b0;
			end
		//For normal case:inside residual_state	
		// 1.entry
		else if (slice_data_state == `residual && residual_state == `rst_residual && !mb_type_general[3])
			trigger_blk4x4_inter_pred <= 1'b1;
		// 2.end of normal
		else if (end_of_one_blk4x4_sum && blk4x4_rec_counter != 23 && !mb_type_general[3])
			trigger_blk4x4_inter_pred <= 1'b1;
		else
			trigger_blk4x4_inter_pred <= 1'b0;
	
	//4. trigger reconstruction sum
	//   Need to align the output of residual(IQIT) and predition(inter/intra)
	wire end_of_one_blk4x4_pred;
	wire end_of_one_blk4x4_res;  //end of one zero or non-zero AC blk4x4 IQIT (NOT DC!)
	reg  blk4x4_res_pred_align;
	
	assign end_of_one_blk4x4_pred = (end_of_one_blk4x4_inter || end_of_one_blk4x4_intra);
	assign end_of_one_blk4x4_res  = (((residual_state == `Intra16x16ACLevel_s || residual_state == `LumaLevel_s || 
								residual_state == `ChromaACLevel_Cb_s || residual_state == `ChromaACLevel_Cr_s) &&  
								(end_of_one_residual_block && TotalCoeff == 0)) || end_of_ACBlk4x4_IQIT)? 1'b1:1'b0; 
	
	//align the completion of prediction and residual decoding
	always @ (posedge clk)
		if (reset_n == 1'b0)
			blk4x4_res_pred_align <= 0;	
		else if (trigger_blk4x4_rec_sum == 1'b1)
			blk4x4_res_pred_align <= 1'b0;
		else if (end_of_one_blk4x4_res && end_of_one_blk4x4_pred) //arrive simultaneously,no align
			blk4x4_res_pred_align <= 1'b0;
		else if (end_of_one_blk4x4_res || end_of_one_blk4x4_pred)
			blk4x4_res_pred_align <= 1'b1;
		
			
	always @ (slice_data_state or residual_state or curr_CBPLuma_IsZero or blk4x4_res_pred_align or 
		end_of_one_blk4x4_pred or end_of_one_blk4x4_res)
		if (slice_data_state == `skip_run_duration)
			trigger_blk4x4_rec_sum <= (end_of_one_blk4x4_pred)? 1'b1:1'b0; 
		// Normal
		else if (residual_state == `Intra16x16ACLevel_s || residual_state == `LumaLevel_s || 
				 residual_state == `ChromaACLevel_Cb_s  || residual_state == `ChromaACLevel_Cr_s)
			begin
				if (curr_CBPLuma_IsZero)
					trigger_blk4x4_rec_sum <= (blk4x4_res_pred_align)? 1'b1:end_of_one_blk4x4_pred;
				else if (end_of_one_blk4x4_res && end_of_one_blk4x4_pred) //arrive simultaneously
					trigger_blk4x4_rec_sum <= 1'b1;
				else if ((end_of_one_blk4x4_res || end_of_one_blk4x4_pred) && blk4x4_res_pred_align)
					trigger_blk4x4_rec_sum <= 1'b1;
				else
					trigger_blk4x4_rec_sum <= 1'b0; 
			end		
		// zero blocks
		else if (residual_state == `Intra16x16ACLevel_0_s || residual_state == `LumaLevel_0_s 
			|| residual_state == `ChromaACLevel_0_s)
			trigger_blk4x4_rec_sum <= (end_of_one_blk4x4_pred || blk4x4_res_pred_align)? 1'b1:1'b0;
		else
			trigger_blk4x4_rec_sum <= 1'b0;
						
	//5.trigger Deblocking Filter
	//assign trigger_MB_DF = (end_of_MB_DEC == 1'b1 && !disable_DF)? 1'b1:1'b0;

	//always @ (posedge clk)
		//$display(" trigger_blk4x4_rec_sum:= %d ", trigger_blk4x4_rec_sum);//////////////////////////////////////


	
endmodule
		
					
		
