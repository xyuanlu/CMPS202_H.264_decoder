//--------------------------------------------------------------------------------------------------
// Design    : nova
// Author(s) : Ke Xu
// Email	   : eexuke@yahoo.com
// File      : Inter_pred_top.v
// Generated : Oct 28, 2005
// Copyright (C) 2008 Ke Xu                
//-------------------------------------------------------------------------------------------------
// Description 
// Top module of Inter prediction, including
// Inter_pred_pipeline.v 		
// Inter_pred_reg_control.v	
// Inter_pred_sliding_window.v 
// Inter_pred_LPE.v			
// Inter_pred_CPE.v			
//-------------------------------------------------------------------------------------------------

// synopsys translate_off
//`include "timescale.v"
// synopsys translate_on
`include "nova_defines.v"

module Inter_pred_top (clk,gclk_Inter_ref_rf,reset_n,mb_num_h,mb_num_v,trigger_blk4x4_inter_pred,blk4x4_rec_counter,
	mb_type_general_bit3,mv_is16x16,mv_below8x8,mvx_CurrMb0,mvx_CurrMb1,mvx_CurrMb2,mvx_CurrMb3,
	mvy_CurrMb0,mvy_CurrMb1,mvy_CurrMb2,mvy_CurrMb3,ref_frame_RAM_dout,
	
	Inter_pred_out0,Inter_pred_out1,Inter_pred_out2,Inter_pred_out3,
	blk4x4_inter_preload_counter,blk4x4_inter_calculate_counter,Inter_chroma2x2_counter,
	mv_below8x8_curr,pos_FracL,end_of_one_blk4x4_inter,Inter_blk4x4_pred_output_valid,
	ref_frame_RAM_rd,ref_frame_RAM_rd_addr);
	input clk;
	input gclk_Inter_ref_rf;
	input reset_n;
	input [3:0] mb_num_h,mb_num_v;
	input trigger_blk4x4_inter_pred;
	input [4:0] blk4x4_rec_counter;
	input mb_type_general_bit3;
	input mv_is16x16;
	input [3:0] mv_below8x8;
	input [31:0] mvx_CurrMb0,mvx_CurrMb1,mvx_CurrMb2,mvx_CurrMb3;
	input [31:0] mvy_CurrMb0,mvy_CurrMb1,mvy_CurrMb2,mvy_CurrMb3;
	input [31:0] ref_frame_RAM_dout;
	
	output [7:0] Inter_pred_out0,Inter_pred_out1,Inter_pred_out2,Inter_pred_out3;
	output [5:0] blk4x4_inter_preload_counter;
	output [3:0] blk4x4_inter_calculate_counter;
	output [1:0] Inter_chroma2x2_counter;
	output mv_below8x8_curr;
	output [3:0] pos_FracL;
	output end_of_one_blk4x4_inter;
	output [1:0] Inter_blk4x4_pred_output_valid;
	output ref_frame_RAM_rd;
	output [13:0] ref_frame_RAM_rd_addr;
	
	wire [7:0] LPE0_out,LPE1_out,LPE2_out,LPE3_out;
	wire [7:0] CPE0_out,CPE1_out,CPE2_out,CPE3_out;
	wire [5:0] blk4x4_inter_preload_counter;
	wire mv_below8x8_curr;
	wire IsInterLuma,IsInterChroma;
	wire Is_InterChromaCopy;
	wire [8:0] xInt_addr_unclip;
	wire [1:0] xInt_org_unclip_1to0;
	wire [2:0] xFracC,yFracC;
	
	wire [7:0] Inter_ref_00_00,Inter_ref_01_00,Inter_ref_02_00,Inter_ref_03_00,Inter_ref_04_00,Inter_ref_05_00;
	wire [7:0] Inter_ref_06_00,Inter_ref_07_00,Inter_ref_08_00,Inter_ref_09_00,Inter_ref_10_00,Inter_ref_11_00,Inter_ref_12_00;
	wire [7:0] Inter_ref_00_01,Inter_ref_01_01,Inter_ref_02_01,Inter_ref_03_01,Inter_ref_04_01,Inter_ref_05_01;
	wire [7:0] Inter_ref_06_01,Inter_ref_07_01,Inter_ref_08_01,Inter_ref_09_01,Inter_ref_10_01,Inter_ref_11_01,Inter_ref_12_01;
	wire [7:0] Inter_ref_00_02,Inter_ref_01_02,Inter_ref_02_02,Inter_ref_03_02,Inter_ref_04_02,Inter_ref_05_02;
	wire [7:0] Inter_ref_06_02,Inter_ref_07_02,Inter_ref_08_02,Inter_ref_09_02,Inter_ref_10_02,Inter_ref_11_02,Inter_ref_12_02;
	wire [7:0] Inter_ref_00_03,Inter_ref_01_03,Inter_ref_02_03,Inter_ref_03_03,Inter_ref_04_03,Inter_ref_05_03;
	wire [7:0] Inter_ref_06_03,Inter_ref_07_03,Inter_ref_08_03,Inter_ref_09_03,Inter_ref_10_03,Inter_ref_11_03,Inter_ref_12_03;
	wire [7:0] Inter_ref_00_04,Inter_ref_01_04,Inter_ref_02_04,Inter_ref_03_04,Inter_ref_04_04,Inter_ref_05_04;
	wire [7:0] Inter_ref_06_04,Inter_ref_07_04,Inter_ref_08_04,Inter_ref_09_04,Inter_ref_10_04,Inter_ref_11_04,Inter_ref_12_04;
	wire [7:0] Inter_ref_00_05,Inter_ref_01_05,Inter_ref_02_05,Inter_ref_03_05,Inter_ref_04_05,Inter_ref_05_05;
	wire [7:0] Inter_ref_06_05,Inter_ref_07_05,Inter_ref_08_05,Inter_ref_09_05,Inter_ref_10_05,Inter_ref_11_05,Inter_ref_12_05;
	wire [7:0] Inter_ref_00_06,Inter_ref_01_06,Inter_ref_02_06,Inter_ref_03_06,Inter_ref_04_06,Inter_ref_05_06;
	wire [7:0] Inter_ref_06_06,Inter_ref_07_06,Inter_ref_08_06,Inter_ref_09_06,Inter_ref_10_06,Inter_ref_11_06,Inter_ref_12_06;
	wire [7:0] Inter_ref_00_07,Inter_ref_01_07,Inter_ref_02_07,Inter_ref_03_07,Inter_ref_04_07,Inter_ref_05_07;
	wire [7:0] Inter_ref_06_07,Inter_ref_07_07,Inter_ref_08_07,Inter_ref_09_07,Inter_ref_10_07,Inter_ref_11_07,Inter_ref_12_07;
	wire [7:0] Inter_ref_00_08,Inter_ref_01_08,Inter_ref_02_08,Inter_ref_03_08,Inter_ref_04_08,Inter_ref_05_08;
	wire [7:0] Inter_ref_06_08,Inter_ref_07_08,Inter_ref_08_08,Inter_ref_09_08,Inter_ref_10_08,Inter_ref_11_08,Inter_ref_12_08;
	wire [7:0] Inter_ref_00_09,Inter_ref_01_09,Inter_ref_02_09,Inter_ref_03_09,Inter_ref_04_09,Inter_ref_05_09;
	wire [7:0] Inter_ref_06_09,Inter_ref_07_09,Inter_ref_08_09,Inter_ref_09_09,Inter_ref_10_09,Inter_ref_11_09,Inter_ref_12_09;
	wire [7:0] Inter_ref_00_10,Inter_ref_01_10,Inter_ref_02_10,Inter_ref_03_10,Inter_ref_04_10,Inter_ref_05_10;
	wire [7:0] Inter_ref_06_10,Inter_ref_07_10,Inter_ref_08_10,Inter_ref_09_10,Inter_ref_10_10,Inter_ref_11_10,Inter_ref_12_10;
	wire [7:0] Inter_ref_00_11,Inter_ref_01_11,Inter_ref_02_11,Inter_ref_03_11,Inter_ref_04_11,Inter_ref_05_11;
	wire [7:0] Inter_ref_06_11,Inter_ref_07_11,Inter_ref_08_11,Inter_ref_09_11,Inter_ref_10_11,Inter_ref_11_11,Inter_ref_12_11;
	wire [7:0] Inter_ref_00_12,Inter_ref_01_12,Inter_ref_02_12,Inter_ref_03_12,Inter_ref_04_12,Inter_ref_05_12;
	wire [7:0] Inter_ref_06_12,Inter_ref_07_12,Inter_ref_08_12,Inter_ref_09_12,Inter_ref_10_12,Inter_ref_11_12,Inter_ref_12_12; 
	
	wire [7:0] Inter_pix_copy0,Inter_pix_copy1,Inter_pix_copy2,Inter_pix_copy3;
	wire [7:0] Inter_H_window_0_0,Inter_H_window_1_0,Inter_H_window_2_0,Inter_H_window_3_0,Inter_H_window_4_0,Inter_H_window_5_0;
	wire [7:0] Inter_H_window_0_1,Inter_H_window_1_1,Inter_H_window_2_1,Inter_H_window_3_1,Inter_H_window_4_1,Inter_H_window_5_1;
	wire [7:0] Inter_H_window_0_2,Inter_H_window_1_2,Inter_H_window_2_2,Inter_H_window_3_2,Inter_H_window_4_2,Inter_H_window_5_2;
	wire [7:0] Inter_H_window_0_3,Inter_H_window_1_3,Inter_H_window_2_3,Inter_H_window_3_3,Inter_H_window_4_3,Inter_H_window_5_3;
	wire [7:0] Inter_H_window_0_4,Inter_H_window_1_4,Inter_H_window_2_4,Inter_H_window_3_4,Inter_H_window_4_4,Inter_H_window_5_4;
	wire [7:0] Inter_H_window_0_5,Inter_H_window_1_5,Inter_H_window_2_5,Inter_H_window_3_5,Inter_H_window_4_5,Inter_H_window_5_5;
	wire [7:0] Inter_H_window_0_6,Inter_H_window_1_6,Inter_H_window_2_6,Inter_H_window_3_6,Inter_H_window_4_6,Inter_H_window_5_6;
	wire [7:0] Inter_H_window_0_7,Inter_H_window_1_7,Inter_H_window_2_7,Inter_H_window_3_7,Inter_H_window_4_7,Inter_H_window_5_7;
	wire [7:0] Inter_H_window_0_8,Inter_H_window_1_8,Inter_H_window_2_8,Inter_H_window_3_8,Inter_H_window_4_8,Inter_H_window_5_8;
	wire [7:0] Inter_V_window_0,Inter_V_window_1,Inter_V_window_2,Inter_V_window_3,Inter_V_window_4;
	wire [7:0] Inter_V_window_5,Inter_V_window_6,Inter_V_window_7,Inter_V_window_8;
	wire [7:0] Inter_C_window_0_0,Inter_C_window_1_0,Inter_C_window_2_0;
	wire [7:0] Inter_C_window_0_1,Inter_C_window_1_1,Inter_C_window_2_1;
	wire [7:0] Inter_C_window_0_2,Inter_C_window_1_2,Inter_C_window_2_2;
	wire [7:0] Inter_bi_window_0,Inter_bi_window_1,Inter_bi_window_2,Inter_bi_window_3;
	
	Inter_pred_pipeline Inter_pred_pipeline(
		.clk(clk),
		.reset_n(reset_n),
		.mb_num_h(mb_num_h),
		.mb_num_v(mb_num_v),
		.trigger_blk4x4_inter_pred(trigger_blk4x4_inter_pred),
		.blk4x4_rec_counter(blk4x4_rec_counter),
		.mb_type_general_bit3(mb_type_general_bit3),
		.mv_is16x16(mv_is16x16),
		.mv_below8x8(mv_below8x8),
		.mvx_CurrMb0(mvx_CurrMb0),
		.mvx_CurrMb1(mvx_CurrMb1),
		.mvx_CurrMb2(mvx_CurrMb2),
		.mvx_CurrMb3(mvx_CurrMb3),
		.mvy_CurrMb0(mvy_CurrMb0),
		.mvy_CurrMb1(mvy_CurrMb1),
		.mvy_CurrMb2(mvy_CurrMb2),
		.mvy_CurrMb3(mvy_CurrMb3),
		.Inter_pix_copy0(Inter_pix_copy0),
		.Inter_pix_copy1(Inter_pix_copy1),
		.Inter_pix_copy2(Inter_pix_copy2),
		.Inter_pix_copy3(Inter_pix_copy3),
		.LPE0_out(LPE0_out),
		.LPE1_out(LPE1_out),
		.LPE2_out(LPE2_out),
		.LPE3_out(LPE3_out),
		.CPE0_out(CPE0_out),
		.CPE1_out(CPE1_out),
		.CPE2_out(CPE2_out),
		.CPE3_out(CPE3_out),
		
		.mv_below8x8_curr(mv_below8x8_curr),
		.blk4x4_inter_preload_counter(blk4x4_inter_preload_counter),
		.blk4x4_inter_calculate_counter(blk4x4_inter_calculate_counter),
		.Inter_chroma2x2_counter(Inter_chroma2x2_counter),
		.end_of_one_blk4x4_inter(end_of_one_blk4x4_inter),
		.IsInterLuma(IsInterLuma),
		.IsInterChroma(IsInterChroma),
		.Is_InterChromaCopy(Is_InterChromaCopy),
		.xInt_addr_unclip(xInt_addr_unclip),
		.xInt_org_unclip_1to0(xInt_org_unclip_1to0),
		.pos_FracL(pos_FracL),
		.xFracC(xFracC),
		.yFracC(yFracC),
		.Inter_pred_out0(Inter_pred_out0),
		.Inter_pred_out1(Inter_pred_out1),
		.Inter_pred_out2(Inter_pred_out2),
		.Inter_pred_out3(Inter_pred_out3),
		.Inter_blk4x4_pred_output_valid(Inter_blk4x4_pred_output_valid),
		.ref_frame_RAM_rd(ref_frame_RAM_rd),
		.ref_frame_RAM_rd_addr(ref_frame_RAM_rd_addr)
		);
	
	Inter_pred_reg_ctrl Inter_pred_reg_ctrl (
		.gclk_Inter_ref_rf(gclk_Inter_ref_rf),
		.reset_n(reset_n),
		.blk4x4_inter_preload_counter(blk4x4_inter_preload_counter),
		.ref_frame_RAM_dout(ref_frame_RAM_dout),
		.IsInterLuma(IsInterLuma),
		.IsInterChroma(IsInterChroma),
		.xInt_addr_unclip(xInt_addr_unclip),
		.xInt_org_unclip_1to0(xInt_org_unclip_1to0),
		.pos_FracL(pos_FracL),
		.xFracC(xFracC),
		.yFracC(yFracC),
		.mv_below8x8_curr(mv_below8x8_curr),
		
		.Inter_ref_00_00(Inter_ref_00_00),
		.Inter_ref_01_00(Inter_ref_01_00),
		.Inter_ref_02_00(Inter_ref_02_00),
		.Inter_ref_03_00(Inter_ref_03_00),
		.Inter_ref_04_00(Inter_ref_04_00),
		.Inter_ref_05_00(Inter_ref_05_00),
		.Inter_ref_06_00(Inter_ref_06_00),
		.Inter_ref_07_00(Inter_ref_07_00),
		.Inter_ref_08_00(Inter_ref_08_00),
		.Inter_ref_09_00(Inter_ref_09_00),
		.Inter_ref_10_00(Inter_ref_10_00),
		.Inter_ref_11_00(Inter_ref_11_00),
		.Inter_ref_12_00(Inter_ref_12_00),
		.Inter_ref_00_01(Inter_ref_00_01),
		.Inter_ref_01_01(Inter_ref_01_01),
		.Inter_ref_02_01(Inter_ref_02_01),
		.Inter_ref_03_01(Inter_ref_03_01),
		.Inter_ref_04_01(Inter_ref_04_01),
		.Inter_ref_05_01(Inter_ref_05_01),
		.Inter_ref_06_01(Inter_ref_06_01),
		.Inter_ref_07_01(Inter_ref_07_01),
		.Inter_ref_08_01(Inter_ref_08_01),
		.Inter_ref_09_01(Inter_ref_09_01),
		.Inter_ref_10_01(Inter_ref_10_01),
		.Inter_ref_11_01(Inter_ref_11_01),
		.Inter_ref_12_01(Inter_ref_12_01),
		.Inter_ref_00_02(Inter_ref_00_02),
		.Inter_ref_01_02(Inter_ref_01_02),
		.Inter_ref_02_02(Inter_ref_02_02),
		.Inter_ref_03_02(Inter_ref_03_02),
		.Inter_ref_04_02(Inter_ref_04_02),
		.Inter_ref_05_02(Inter_ref_05_02),
		.Inter_ref_06_02(Inter_ref_06_02),
		.Inter_ref_07_02(Inter_ref_07_02),
		.Inter_ref_08_02(Inter_ref_08_02),
		.Inter_ref_09_02(Inter_ref_09_02),
		.Inter_ref_10_02(Inter_ref_10_02),
		.Inter_ref_11_02(Inter_ref_11_02),
		.Inter_ref_12_02(Inter_ref_12_02),
		.Inter_ref_00_03(Inter_ref_00_03),
		.Inter_ref_01_03(Inter_ref_01_03),
		.Inter_ref_02_03(Inter_ref_02_03),
		.Inter_ref_03_03(Inter_ref_03_03),
		.Inter_ref_04_03(Inter_ref_04_03),
		.Inter_ref_05_03(Inter_ref_05_03),
		.Inter_ref_06_03(Inter_ref_06_03),
		.Inter_ref_07_03(Inter_ref_07_03),
		.Inter_ref_08_03(Inter_ref_08_03),
		.Inter_ref_09_03(Inter_ref_09_03),
		.Inter_ref_10_03(Inter_ref_10_03),
		.Inter_ref_11_03(Inter_ref_11_03),
		.Inter_ref_12_03(Inter_ref_12_03),
		.Inter_ref_00_04(Inter_ref_00_04),
		.Inter_ref_01_04(Inter_ref_01_04),
		.Inter_ref_02_04(Inter_ref_02_04),
		.Inter_ref_03_04(Inter_ref_03_04),
		.Inter_ref_04_04(Inter_ref_04_04),
		.Inter_ref_05_04(Inter_ref_05_04),
		.Inter_ref_06_04(Inter_ref_06_04),
		.Inter_ref_07_04(Inter_ref_07_04),
		.Inter_ref_08_04(Inter_ref_08_04),
		.Inter_ref_09_04(Inter_ref_09_04),
		.Inter_ref_10_04(Inter_ref_10_04),
		.Inter_ref_11_04(Inter_ref_11_04),
		.Inter_ref_12_04(Inter_ref_12_04),
		.Inter_ref_00_05(Inter_ref_00_05),
		.Inter_ref_01_05(Inter_ref_01_05),
		.Inter_ref_02_05(Inter_ref_02_05),
		.Inter_ref_03_05(Inter_ref_03_05),
		.Inter_ref_04_05(Inter_ref_04_05),
		.Inter_ref_05_05(Inter_ref_05_05),
		.Inter_ref_06_05(Inter_ref_06_05),
		.Inter_ref_07_05(Inter_ref_07_05),
		.Inter_ref_08_05(Inter_ref_08_05),
		.Inter_ref_09_05(Inter_ref_09_05),
		.Inter_ref_10_05(Inter_ref_10_05),
		.Inter_ref_11_05(Inter_ref_11_05),
		.Inter_ref_12_05(Inter_ref_12_05),
		.Inter_ref_00_06(Inter_ref_00_06),
		.Inter_ref_01_06(Inter_ref_01_06),
		.Inter_ref_02_06(Inter_ref_02_06),
		.Inter_ref_03_06(Inter_ref_03_06),
		.Inter_ref_04_06(Inter_ref_04_06),
		.Inter_ref_05_06(Inter_ref_05_06),
		.Inter_ref_06_06(Inter_ref_06_06),
		.Inter_ref_07_06(Inter_ref_07_06),
		.Inter_ref_08_06(Inter_ref_08_06),
		.Inter_ref_09_06(Inter_ref_09_06),
		.Inter_ref_10_06(Inter_ref_10_06),
		.Inter_ref_11_06(Inter_ref_11_06),
		.Inter_ref_12_06(Inter_ref_12_06),
		.Inter_ref_00_07(Inter_ref_00_07),
		.Inter_ref_01_07(Inter_ref_01_07),
		.Inter_ref_02_07(Inter_ref_02_07),
		.Inter_ref_03_07(Inter_ref_03_07),
		.Inter_ref_04_07(Inter_ref_04_07),
		.Inter_ref_05_07(Inter_ref_05_07),
		.Inter_ref_06_07(Inter_ref_06_07),
		.Inter_ref_07_07(Inter_ref_07_07),
		.Inter_ref_08_07(Inter_ref_08_07),
		.Inter_ref_09_07(Inter_ref_09_07),
		.Inter_ref_10_07(Inter_ref_10_07),
		.Inter_ref_11_07(Inter_ref_11_07),
		.Inter_ref_12_07(Inter_ref_12_07),
		.Inter_ref_00_08(Inter_ref_00_08),
		.Inter_ref_01_08(Inter_ref_01_08),
		.Inter_ref_02_08(Inter_ref_02_08),
		.Inter_ref_03_08(Inter_ref_03_08),
		.Inter_ref_04_08(Inter_ref_04_08),
		.Inter_ref_05_08(Inter_ref_05_08),
		.Inter_ref_06_08(Inter_ref_06_08),
		.Inter_ref_07_08(Inter_ref_07_08),
		.Inter_ref_08_08(Inter_ref_08_08),
		.Inter_ref_09_08(Inter_ref_09_08),
		.Inter_ref_10_08(Inter_ref_10_08),
		.Inter_ref_11_08(Inter_ref_11_08),
		.Inter_ref_12_08(Inter_ref_12_08),
		.Inter_ref_00_09(Inter_ref_00_09),
		.Inter_ref_01_09(Inter_ref_01_09),
		.Inter_ref_02_09(Inter_ref_02_09),
		.Inter_ref_03_09(Inter_ref_03_09),
		.Inter_ref_04_09(Inter_ref_04_09),
		.Inter_ref_05_09(Inter_ref_05_09),
		.Inter_ref_06_09(Inter_ref_06_09),
		.Inter_ref_07_09(Inter_ref_07_09),
		.Inter_ref_08_09(Inter_ref_08_09),
		.Inter_ref_09_09(Inter_ref_09_09),
		.Inter_ref_10_09(Inter_ref_10_09),
		.Inter_ref_11_09(Inter_ref_11_09),
		.Inter_ref_12_09(Inter_ref_12_09),
		.Inter_ref_00_10(Inter_ref_00_10),
		.Inter_ref_01_10(Inter_ref_01_10),
		.Inter_ref_02_10(Inter_ref_02_10),
		.Inter_ref_03_10(Inter_ref_03_10),
		.Inter_ref_04_10(Inter_ref_04_10),
		.Inter_ref_05_10(Inter_ref_05_10),
		.Inter_ref_06_10(Inter_ref_06_10),
		.Inter_ref_07_10(Inter_ref_07_10),
		.Inter_ref_08_10(Inter_ref_08_10),
		.Inter_ref_09_10(Inter_ref_09_10),
		.Inter_ref_10_10(Inter_ref_10_10),
		.Inter_ref_11_10(Inter_ref_11_10),
		.Inter_ref_12_10(Inter_ref_12_10),
		.Inter_ref_00_11(Inter_ref_00_11),
		.Inter_ref_01_11(Inter_ref_01_11),
		.Inter_ref_02_11(Inter_ref_02_11),
		.Inter_ref_03_11(Inter_ref_03_11),
		.Inter_ref_04_11(Inter_ref_04_11),
		.Inter_ref_05_11(Inter_ref_05_11),
		.Inter_ref_06_11(Inter_ref_06_11),
		.Inter_ref_07_11(Inter_ref_07_11),
		.Inter_ref_08_11(Inter_ref_08_11),
		.Inter_ref_09_11(Inter_ref_09_11),
		.Inter_ref_10_11(Inter_ref_10_11),
		.Inter_ref_11_11(Inter_ref_11_11),
		.Inter_ref_12_11(Inter_ref_12_11),
		.Inter_ref_00_12(Inter_ref_00_12),
		.Inter_ref_01_12(Inter_ref_01_12),
		.Inter_ref_02_12(Inter_ref_02_12),
		.Inter_ref_03_12(Inter_ref_03_12),
		.Inter_ref_04_12(Inter_ref_04_12),
		.Inter_ref_05_12(Inter_ref_05_12),
		.Inter_ref_06_12(Inter_ref_06_12),
		.Inter_ref_07_12(Inter_ref_07_12),
		.Inter_ref_08_12(Inter_ref_08_12),
		.Inter_ref_09_12(Inter_ref_09_12),
		.Inter_ref_10_12(Inter_ref_10_12),
		.Inter_ref_11_12(Inter_ref_11_12),
		.Inter_ref_12_12(Inter_ref_12_12)
		);
	Inter_pred_sliding_window Inter_pred_sliding_window (
		.IsInterLuma(IsInterLuma),
		.IsInterChroma(IsInterChroma),
		.Is_InterChromaCopy(Is_InterChromaCopy),
		.mv_below8x8_curr(mv_below8x8_curr),
		.pos_FracL(pos_FracL),
		.blk4x4_rec_counter_1to0(blk4x4_rec_counter[1:0]),
		.blk4x4_inter_calculate_counter(blk4x4_inter_calculate_counter),
	 	.Inter_ref_00_00(Inter_ref_00_00),
		.Inter_ref_01_00(Inter_ref_01_00),
		.Inter_ref_02_00(Inter_ref_02_00),
		.Inter_ref_03_00(Inter_ref_03_00),
		.Inter_ref_04_00(Inter_ref_04_00),
		.Inter_ref_05_00(Inter_ref_05_00),
		.Inter_ref_06_00(Inter_ref_06_00),
		.Inter_ref_07_00(Inter_ref_07_00),
		.Inter_ref_08_00(Inter_ref_08_00),
		.Inter_ref_09_00(Inter_ref_09_00),
		.Inter_ref_10_00(Inter_ref_10_00),
		.Inter_ref_11_00(Inter_ref_11_00),
		.Inter_ref_12_00(Inter_ref_12_00),
		.Inter_ref_00_01(Inter_ref_00_01),
		.Inter_ref_01_01(Inter_ref_01_01),
		.Inter_ref_02_01(Inter_ref_02_01),
		.Inter_ref_03_01(Inter_ref_03_01),
		.Inter_ref_04_01(Inter_ref_04_01),
		.Inter_ref_05_01(Inter_ref_05_01),
		.Inter_ref_06_01(Inter_ref_06_01),
		.Inter_ref_07_01(Inter_ref_07_01),
		.Inter_ref_08_01(Inter_ref_08_01),
		.Inter_ref_09_01(Inter_ref_09_01),
		.Inter_ref_10_01(Inter_ref_10_01),
		.Inter_ref_11_01(Inter_ref_11_01),
		.Inter_ref_12_01(Inter_ref_12_01),
		.Inter_ref_00_02(Inter_ref_00_02),
		.Inter_ref_01_02(Inter_ref_01_02),
		.Inter_ref_02_02(Inter_ref_02_02),
		.Inter_ref_03_02(Inter_ref_03_02),
		.Inter_ref_04_02(Inter_ref_04_02),
		.Inter_ref_05_02(Inter_ref_05_02),
		.Inter_ref_06_02(Inter_ref_06_02),
		.Inter_ref_07_02(Inter_ref_07_02),
		.Inter_ref_08_02(Inter_ref_08_02),
		.Inter_ref_09_02(Inter_ref_09_02),
		.Inter_ref_10_02(Inter_ref_10_02),
		.Inter_ref_11_02(Inter_ref_11_02),
		.Inter_ref_12_02(Inter_ref_12_02),
		.Inter_ref_00_03(Inter_ref_00_03),
		.Inter_ref_01_03(Inter_ref_01_03),
		.Inter_ref_02_03(Inter_ref_02_03),
		.Inter_ref_03_03(Inter_ref_03_03),
		.Inter_ref_04_03(Inter_ref_04_03),
		.Inter_ref_05_03(Inter_ref_05_03),
		.Inter_ref_06_03(Inter_ref_06_03),
		.Inter_ref_07_03(Inter_ref_07_03),
		.Inter_ref_08_03(Inter_ref_08_03),
		.Inter_ref_09_03(Inter_ref_09_03),
		.Inter_ref_10_03(Inter_ref_10_03),
		.Inter_ref_11_03(Inter_ref_11_03),
		.Inter_ref_12_03(Inter_ref_12_03),
		.Inter_ref_00_04(Inter_ref_00_04),
		.Inter_ref_01_04(Inter_ref_01_04),
		.Inter_ref_02_04(Inter_ref_02_04),
		.Inter_ref_03_04(Inter_ref_03_04),
		.Inter_ref_04_04(Inter_ref_04_04),
		.Inter_ref_05_04(Inter_ref_05_04),
		.Inter_ref_06_04(Inter_ref_06_04),
		.Inter_ref_07_04(Inter_ref_07_04),
		.Inter_ref_08_04(Inter_ref_08_04),
		.Inter_ref_09_04(Inter_ref_09_04),
		.Inter_ref_10_04(Inter_ref_10_04),
		.Inter_ref_11_04(Inter_ref_11_04),
		.Inter_ref_12_04(Inter_ref_12_04),
		.Inter_ref_00_05(Inter_ref_00_05),
		.Inter_ref_01_05(Inter_ref_01_05),
		.Inter_ref_02_05(Inter_ref_02_05),
		.Inter_ref_03_05(Inter_ref_03_05),
		.Inter_ref_04_05(Inter_ref_04_05),
		.Inter_ref_05_05(Inter_ref_05_05),
		.Inter_ref_06_05(Inter_ref_06_05),
		.Inter_ref_07_05(Inter_ref_07_05),
		.Inter_ref_08_05(Inter_ref_08_05),
		.Inter_ref_09_05(Inter_ref_09_05),
		.Inter_ref_10_05(Inter_ref_10_05),
		.Inter_ref_11_05(Inter_ref_11_05),
		.Inter_ref_12_05(Inter_ref_12_05),
		.Inter_ref_00_06(Inter_ref_00_06),
		.Inter_ref_01_06(Inter_ref_01_06),
		.Inter_ref_02_06(Inter_ref_02_06),
		.Inter_ref_03_06(Inter_ref_03_06),
		.Inter_ref_04_06(Inter_ref_04_06),
		.Inter_ref_05_06(Inter_ref_05_06),
		.Inter_ref_06_06(Inter_ref_06_06),
		.Inter_ref_07_06(Inter_ref_07_06),
		.Inter_ref_08_06(Inter_ref_08_06),
		.Inter_ref_09_06(Inter_ref_09_06),
		.Inter_ref_10_06(Inter_ref_10_06),
		.Inter_ref_11_06(Inter_ref_11_06),
		.Inter_ref_12_06(Inter_ref_12_06),
		.Inter_ref_00_07(Inter_ref_00_07),
		.Inter_ref_01_07(Inter_ref_01_07),
		.Inter_ref_02_07(Inter_ref_02_07),
		.Inter_ref_03_07(Inter_ref_03_07),
		.Inter_ref_04_07(Inter_ref_04_07),
		.Inter_ref_05_07(Inter_ref_05_07),
		.Inter_ref_06_07(Inter_ref_06_07),
		.Inter_ref_07_07(Inter_ref_07_07),
		.Inter_ref_08_07(Inter_ref_08_07),
		.Inter_ref_09_07(Inter_ref_09_07),
		.Inter_ref_10_07(Inter_ref_10_07),
		.Inter_ref_11_07(Inter_ref_11_07),
		.Inter_ref_12_07(Inter_ref_12_07),
		.Inter_ref_00_08(Inter_ref_00_08),
		.Inter_ref_01_08(Inter_ref_01_08),
		.Inter_ref_02_08(Inter_ref_02_08),
		.Inter_ref_03_08(Inter_ref_03_08),
		.Inter_ref_04_08(Inter_ref_04_08),
		.Inter_ref_05_08(Inter_ref_05_08),
		.Inter_ref_06_08(Inter_ref_06_08),
		.Inter_ref_07_08(Inter_ref_07_08),
		.Inter_ref_08_08(Inter_ref_08_08),
		.Inter_ref_09_08(Inter_ref_09_08),
		.Inter_ref_10_08(Inter_ref_10_08),
		.Inter_ref_11_08(Inter_ref_11_08),
		.Inter_ref_12_08(Inter_ref_12_08),
		.Inter_ref_00_09(Inter_ref_00_09),
		.Inter_ref_01_09(Inter_ref_01_09),
		.Inter_ref_02_09(Inter_ref_02_09),
		.Inter_ref_03_09(Inter_ref_03_09),
		.Inter_ref_04_09(Inter_ref_04_09),
		.Inter_ref_05_09(Inter_ref_05_09),
		.Inter_ref_06_09(Inter_ref_06_09),
		.Inter_ref_07_09(Inter_ref_07_09),
		.Inter_ref_08_09(Inter_ref_08_09),
		.Inter_ref_09_09(Inter_ref_09_09),
		.Inter_ref_10_09(Inter_ref_10_09),
		.Inter_ref_11_09(Inter_ref_11_09),
		.Inter_ref_12_09(Inter_ref_12_09),
		.Inter_ref_00_10(Inter_ref_00_10),
		.Inter_ref_01_10(Inter_ref_01_10),
		.Inter_ref_02_10(Inter_ref_02_10),
		.Inter_ref_03_10(Inter_ref_03_10),
		.Inter_ref_04_10(Inter_ref_04_10),
		.Inter_ref_05_10(Inter_ref_05_10),
		.Inter_ref_06_10(Inter_ref_06_10),
		.Inter_ref_07_10(Inter_ref_07_10),
		.Inter_ref_08_10(Inter_ref_08_10),
		.Inter_ref_09_10(Inter_ref_09_10),
		.Inter_ref_10_10(Inter_ref_10_10),
		.Inter_ref_11_10(Inter_ref_11_10),
		.Inter_ref_12_10(Inter_ref_12_10),
		.Inter_ref_00_11(Inter_ref_00_11),
		.Inter_ref_01_11(Inter_ref_01_11),
		.Inter_ref_02_11(Inter_ref_02_11),
		.Inter_ref_03_11(Inter_ref_03_11),
		.Inter_ref_04_11(Inter_ref_04_11),
		.Inter_ref_05_11(Inter_ref_05_11),
		.Inter_ref_06_11(Inter_ref_06_11),
		.Inter_ref_07_11(Inter_ref_07_11),
		.Inter_ref_08_11(Inter_ref_08_11),
		.Inter_ref_09_11(Inter_ref_09_11),
		.Inter_ref_10_11(Inter_ref_10_11),
		.Inter_ref_11_11(Inter_ref_11_11),
		.Inter_ref_12_11(Inter_ref_12_11),
		.Inter_ref_00_12(Inter_ref_00_12),
		.Inter_ref_01_12(Inter_ref_01_12),
		.Inter_ref_02_12(Inter_ref_02_12),
		.Inter_ref_03_12(Inter_ref_03_12),
		.Inter_ref_04_12(Inter_ref_04_12),
		.Inter_ref_05_12(Inter_ref_05_12),
		.Inter_ref_06_12(Inter_ref_06_12),
		.Inter_ref_07_12(Inter_ref_07_12),
		.Inter_ref_08_12(Inter_ref_08_12),
		.Inter_ref_09_12(Inter_ref_09_12),
		.Inter_ref_10_12(Inter_ref_10_12),
		.Inter_ref_11_12(Inter_ref_11_12),
		.Inter_ref_12_12(Inter_ref_12_12),
	
		.Inter_pix_copy0(Inter_pix_copy0),
		.Inter_pix_copy1(Inter_pix_copy1),
		.Inter_pix_copy2(Inter_pix_copy2),
		.Inter_pix_copy3(Inter_pix_copy3),
		.Inter_H_window_0_0(Inter_H_window_0_0),
		.Inter_H_window_1_0(Inter_H_window_1_0),
		.Inter_H_window_2_0(Inter_H_window_2_0),
		.Inter_H_window_3_0(Inter_H_window_3_0),
		.Inter_H_window_4_0(Inter_H_window_4_0),
		.Inter_H_window_5_0(Inter_H_window_5_0),
		.Inter_H_window_0_1(Inter_H_window_0_1),
		.Inter_H_window_1_1(Inter_H_window_1_1),
		.Inter_H_window_2_1(Inter_H_window_2_1),
		.Inter_H_window_3_1(Inter_H_window_3_1),
		.Inter_H_window_4_1(Inter_H_window_4_1),
		.Inter_H_window_5_1(Inter_H_window_5_1),
		.Inter_H_window_0_2(Inter_H_window_0_2),
		.Inter_H_window_1_2(Inter_H_window_1_2),
		.Inter_H_window_2_2(Inter_H_window_2_2),
		.Inter_H_window_3_2(Inter_H_window_3_2),
		.Inter_H_window_4_2(Inter_H_window_4_2),
		.Inter_H_window_5_2(Inter_H_window_5_2),
		.Inter_H_window_0_3(Inter_H_window_0_3),
		.Inter_H_window_1_3(Inter_H_window_1_3),
		.Inter_H_window_2_3(Inter_H_window_2_3),
		.Inter_H_window_3_3(Inter_H_window_3_3),
		.Inter_H_window_4_3(Inter_H_window_4_3),
		.Inter_H_window_5_3(Inter_H_window_5_3),
		.Inter_H_window_0_4(Inter_H_window_0_4),
		.Inter_H_window_1_4(Inter_H_window_1_4),
		.Inter_H_window_2_4(Inter_H_window_2_4),
		.Inter_H_window_3_4(Inter_H_window_3_4),
		.Inter_H_window_4_4(Inter_H_window_4_4),
		.Inter_H_window_5_4(Inter_H_window_5_4),
		.Inter_H_window_0_5(Inter_H_window_0_5),
		.Inter_H_window_1_5(Inter_H_window_1_5),
		.Inter_H_window_2_5(Inter_H_window_2_5),
		.Inter_H_window_3_5(Inter_H_window_3_5),
		.Inter_H_window_4_5(Inter_H_window_4_5),
		.Inter_H_window_5_5(Inter_H_window_5_5),
		.Inter_H_window_0_6(Inter_H_window_0_6),
		.Inter_H_window_1_6(Inter_H_window_1_6),
		.Inter_H_window_2_6(Inter_H_window_2_6),
		.Inter_H_window_3_6(Inter_H_window_3_6),
		.Inter_H_window_4_6(Inter_H_window_4_6),
		.Inter_H_window_5_6(Inter_H_window_5_6),
		.Inter_H_window_0_7(Inter_H_window_0_7),
		.Inter_H_window_1_7(Inter_H_window_1_7),
		.Inter_H_window_2_7(Inter_H_window_2_7),
		.Inter_H_window_3_7(Inter_H_window_3_7),
		.Inter_H_window_4_7(Inter_H_window_4_7),
		.Inter_H_window_5_7(Inter_H_window_5_7),
		.Inter_H_window_0_8(Inter_H_window_0_8),
		.Inter_H_window_1_8(Inter_H_window_1_8),
		.Inter_H_window_2_8(Inter_H_window_2_8),
		.Inter_H_window_3_8(Inter_H_window_3_8),
		.Inter_H_window_4_8(Inter_H_window_4_8),
		.Inter_H_window_5_8(Inter_H_window_5_8),
		.Inter_V_window_0(Inter_V_window_0), 
		.Inter_V_window_1(Inter_V_window_1), 
		.Inter_V_window_2(Inter_V_window_2), 
		.Inter_V_window_3(Inter_V_window_3), 
		.Inter_V_window_4(Inter_V_window_4), 
		.Inter_V_window_5(Inter_V_window_5), 
		.Inter_V_window_6(Inter_V_window_6),
		.Inter_V_window_7(Inter_V_window_7),
		.Inter_V_window_8(Inter_V_window_8),
		.Inter_C_window_0_0(Inter_C_window_0_0),
		.Inter_C_window_1_0(Inter_C_window_1_0),
		.Inter_C_window_2_0(Inter_C_window_2_0),
		.Inter_C_window_0_1(Inter_C_window_0_1),
		.Inter_C_window_1_1(Inter_C_window_1_1),
		.Inter_C_window_2_1(Inter_C_window_2_1),
		.Inter_C_window_0_2(Inter_C_window_0_2),
		.Inter_C_window_1_2(Inter_C_window_1_2),
		.Inter_C_window_2_2(Inter_C_window_2_2),
		.Inter_bi_window_0(Inter_bi_window_0),
		.Inter_bi_window_1(Inter_bi_window_1),
		.Inter_bi_window_2(Inter_bi_window_2),
		.Inter_bi_window_3(Inter_bi_window_3)
		);
	                        
	Inter_pred_LPE Inter_pred_LPE (
		.clk(clk),      
		.reset_n(reset_n),
		.pos_FracL(pos_FracL),
		.IsInterLuma(IsInterLuma),
		.blk4x4_inter_calculate_counter(blk4x4_inter_calculate_counter),
		.Inter_H_window_0_0(Inter_H_window_0_0),
		.Inter_H_window_1_0(Inter_H_window_1_0),
		.Inter_H_window_2_0(Inter_H_window_2_0),
		.Inter_H_window_3_0(Inter_H_window_3_0),
		.Inter_H_window_4_0(Inter_H_window_4_0),
		.Inter_H_window_5_0(Inter_H_window_5_0),
		.Inter_H_window_0_1(Inter_H_window_0_1),
		.Inter_H_window_1_1(Inter_H_window_1_1),
		.Inter_H_window_2_1(Inter_H_window_2_1),
		.Inter_H_window_3_1(Inter_H_window_3_1),
		.Inter_H_window_4_1(Inter_H_window_4_1),
		.Inter_H_window_5_1(Inter_H_window_5_1),
		.Inter_H_window_0_2(Inter_H_window_0_2),
		.Inter_H_window_1_2(Inter_H_window_1_2),
		.Inter_H_window_2_2(Inter_H_window_2_2),
		.Inter_H_window_3_2(Inter_H_window_3_2),
		.Inter_H_window_4_2(Inter_H_window_4_2),
		.Inter_H_window_5_2(Inter_H_window_5_2),
		.Inter_H_window_0_3(Inter_H_window_0_3),
		.Inter_H_window_1_3(Inter_H_window_1_3),
		.Inter_H_window_2_3(Inter_H_window_2_3),
		.Inter_H_window_3_3(Inter_H_window_3_3),
		.Inter_H_window_4_3(Inter_H_window_4_3),
		.Inter_H_window_5_3(Inter_H_window_5_3),
		.Inter_H_window_0_4(Inter_H_window_0_4),
		.Inter_H_window_1_4(Inter_H_window_1_4),
		.Inter_H_window_2_4(Inter_H_window_2_4),
		.Inter_H_window_3_4(Inter_H_window_3_4),
		.Inter_H_window_4_4(Inter_H_window_4_4),
		.Inter_H_window_5_4(Inter_H_window_5_4),
		.Inter_H_window_0_5(Inter_H_window_0_5),
		.Inter_H_window_1_5(Inter_H_window_1_5),
		.Inter_H_window_2_5(Inter_H_window_2_5),
		.Inter_H_window_3_5(Inter_H_window_3_5),
		.Inter_H_window_4_5(Inter_H_window_4_5),
		.Inter_H_window_5_5(Inter_H_window_5_5),
		.Inter_H_window_0_6(Inter_H_window_0_6),
		.Inter_H_window_1_6(Inter_H_window_1_6),
		.Inter_H_window_2_6(Inter_H_window_2_6),
		.Inter_H_window_3_6(Inter_H_window_3_6),
		.Inter_H_window_4_6(Inter_H_window_4_6),
		.Inter_H_window_5_6(Inter_H_window_5_6),
		.Inter_H_window_0_7(Inter_H_window_0_7),
		.Inter_H_window_1_7(Inter_H_window_1_7),
		.Inter_H_window_2_7(Inter_H_window_2_7),
		.Inter_H_window_3_7(Inter_H_window_3_7),
		.Inter_H_window_4_7(Inter_H_window_4_7),
		.Inter_H_window_5_7(Inter_H_window_5_7),
		.Inter_H_window_0_8(Inter_H_window_0_8),
		.Inter_H_window_1_8(Inter_H_window_1_8),
		.Inter_H_window_2_8(Inter_H_window_2_8),
		.Inter_H_window_3_8(Inter_H_window_3_8),
		.Inter_H_window_4_8(Inter_H_window_4_8),
		.Inter_H_window_5_8(Inter_H_window_5_8),
		.Inter_V_window_0(Inter_V_window_0), 
		.Inter_V_window_1(Inter_V_window_1), 
		.Inter_V_window_2(Inter_V_window_2), 
		.Inter_V_window_3(Inter_V_window_3), 
		.Inter_V_window_4(Inter_V_window_4), 
		.Inter_V_window_5(Inter_V_window_5), 
		.Inter_V_window_6(Inter_V_window_6),
		.Inter_V_window_7(Inter_V_window_7),
		.Inter_V_window_8(Inter_V_window_8),
		.Inter_bi_window_0(Inter_bi_window_0),
		.Inter_bi_window_1(Inter_bi_window_1),
		.Inter_bi_window_2(Inter_bi_window_2),
		.Inter_bi_window_3(Inter_bi_window_3),
	
		.LPE0_out(LPE0_out),
		.LPE1_out(LPE1_out),
		.LPE2_out(LPE2_out),
		.LPE3_out(LPE3_out)
		);
	Inter_pred_CPE Inter_pred_CPE (
		.xFracC(xFracC),
		.yFracC(yFracC),
		.Inter_C_window_0_0(Inter_C_window_0_0),
		.Inter_C_window_1_0(Inter_C_window_1_0),
		.Inter_C_window_2_0(Inter_C_window_2_0),
		.Inter_C_window_0_1(Inter_C_window_0_1),
		.Inter_C_window_1_1(Inter_C_window_1_1),
		.Inter_C_window_2_1(Inter_C_window_2_1),
		.Inter_C_window_0_2(Inter_C_window_0_2),
		.Inter_C_window_1_2(Inter_C_window_1_2),
		.Inter_C_window_2_2(Inter_C_window_2_2),
		.CPE0_out(CPE0_out),
		.CPE1_out(CPE1_out),
		.CPE2_out(CPE2_out),
		.CPE3_out(CPE3_out)
		);
endmodule
	
